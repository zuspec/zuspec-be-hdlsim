module XtorComponent(

);

endmodule
