module CounterControlXtor(
  output logic clk_out,
  output logic rst_out,
  output logic enable_out,
  input logic [7:0] count_in
);

endmodule
